library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_64x8_sync is 
	port (Clock  	: in std_logic;
			Address	: in std_logic_vector(5 downto 0);
			data_out	: out std_logic_vector(7 downto 0));
end entity;

architecture rom_64x8_sync_arch of rom_64x8_sync is

	type ROM_type is array (0 to 63) of std_logic_vector(7 downto 0);
	
	constant ROM : ROM_type := (0  => "00000000",
										 1  => "00010001",
										 2  => "00100010",
										 3  => "00110011",
										 4  => "01000100",
										 5  => "01010101",
										 6  => "01100110",
										 7  => "01110111",
										 8  => "10001000",
										 9  => "10011001",
										 10 => "10101010",
										 11 => "10111011",
										 12 => "11001100",
										 13 => "11011101",
										 14 => "11101110",
										 15 => "11111111",
										 16 => "11111111",
										 17 => "11101110",
										 18 => "11011101",
										 19 => "11001100",
										 20 => "10111011",
										 21 => "10101010",
										 22 => "10011001",
										 23 => "10001000",
										 24 => "01110111",
										 25 => "01100110",
										 26 => "01010101",
										 27 => "01000100",
										 28 => "00110011",
										 29 => "00100010",
										 30 => "00010001",
										 31 => "00000000",
										 32 => "00000000",
										 33 => "00000000",
										 34 => "00000000",
										 35 => "00000000",
										 36 => "00000000",
										 37 => "00000000",
										 38 => "00000000",
										 39 => "00000000",
										 40 => "00000000",
										 41 => "00000000",
										 42 => "00000000",
										 43 => "00000000",
										 44 => "00000000",
										 45 => "00000000",
										 46 => "00000000",
										 47 => "00000000",
										 48 => "00000000",
										 49 => "00000000",
										 50 => "00000000",
										 51 => "00000000",
										 52 => "00000000",
										 53 => "00000000",
										 54 => "00000000",
										 55 => "00000000",
										 56 => "00000000",
										 57 => "00000000",
										 58 => "00000000",
										 59 => "00000000",
										 60 => "00000000",
										 61 => "00000000",
										 62 => "00000000",
										 63 => "00000000");
										 
	
	begin
		MEMORY : process (Clock)
			begin 
				if (rising_edge(Clock)) then
					data_out <= ROM (to_integer(unsigned(address)));
				end if;
		end process;	
		
end architecture;